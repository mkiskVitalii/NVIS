library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity my_mult is
    port(
        DIN  : in  STD_LOGIC_VECTOR(31 downto 0);
        DOUT : out STD_LOGIC_VECTOR(31 downto 0)
    );
end my_mult;

architecture my_mult of my_mult is
    signal X_L1, X_L3, X_L8, X_L9, X_L10, X_L16, X_L17, X_L19, X_L20, X_L21, X_L24, X_L25, X_L27, X_L28, X_L30 : STD_LOGIC_VECTOR(63 downto 0) := (others => '0');
    signal X_L1_L3, X_L8_L9, X_L10_L16, X_L17_L19, X_L20_L21, X_L24_L25, X_L27_L28 : STD_LOGIC_VECTOR(63 downto 0) := (others => '0');
    signal X_L1_L3_L8_L9, X_L10_L16_L17_L19, X_L20_L21_L24_L25, X_L27_L28_L30 : STD_LOGIC_VECTOR(63 downto 0) := (others => '0');
    signal X_L1_L3_L8_L9_L10_L16_L17_19, X_L20_L21_L24_L25_L27_L28_L30 : STD_LOGIC_VECTOR(63 downto 0) := (others => '0');
    signal Y : STD_LOGIC_VECTOR(63 downto 0) := (others => '0');
begin
    X_L1  <= "0000000000000000000000000000000" & DIN & "0";
    X_L3  <= "00000000000000000000000000000" & DIN & "000";
    X_L8  <= "000000000000000000000000" & DIN & "00000000";
    X_L9  <= "00000000000000000000000" & DIN & "000000000";
    X_L10 <= "0000000000000000000000" & DIN & "0000000000";
    X_L16 <= "0000000000000000" & DIN & "0000000000000000";
    X_L17 <= "000000000000000" & DIN & "00000000000000000";
    X_L19 <= "0000000000000" & DIN & "0000000000000000000";
    X_L20 <= "000000000000" & DIN & "00000000000000000000";
    X_L21 <= "00000000000" & DIN & "000000000000000000000";
    X_L24 <= "00000000" & DIN & "000000000000000000000000";
    X_L25 <= "0000000" & DIN & "0000000000000000000000000";
    X_L27 <= "00000" & DIN & "000000000000000000000000000";
    X_L28 <= "0000" & DIN & "0000000000000000000000000000";
    X_L30 <= "00" & DIN & "000000000000000000000000000000";

    X_L1_L3 <= X_L1 + X_L3;
    X_L8_L9 <= X_L8 + X_L9;
    X_L10_L16 <= X_L10 + X_L16;
    X_L17_L19 <= X_L17 + X_L19;
    X_L20_L21 <= X_L20 + X_L21;
    X_L24_L25 <= X_L24 + X_L25;
    X_L27_L28 <= X_L27 + X_L28;

    X_L1_L3_L8_L9 <= X_L1_L3 + X_L8_L9;
    X_L10_L16_L17_L19 <= X_L10_L16 + X_L17_L19;
    X_L20_L21_L24_L25 <= X_L20_L21 + X_L24_L25;
    X_L27_L28_L30 <= X_L27_L28 + X_L30;

    X_L1_L3_L8_L9_L10_L16_L17_19 <= X_L1_L3_L8_L9 + X_L10_L16_L17_L19;
    X_L20_L21_L24_L25_L27_L28_L30 <= X_L20_L21_L24_L25 + X_L27_L28_L30;

    Y <= X_L1_L3_L8_L9_L10_L16_L17_19 + X_L20_L21_L24_L25_L27_L28_L30;
    DOUT <= Y(63 downto 32);
end my_mult;