library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity my_mult is
    port(
        DIN  : in  STD_LOGIC_VECTOR(31 downto 0);
        DOUT : out STD_LOGIC_VECTOR(31 downto 0)
    );
end my_mult;

architecture my_mult of my_mult is
    signal X_L1, X_L3, X_L8, X_L11, X_L16, X_L18, X_L22, X_L24, X_L26, X_L29, X_L30 : STD_LOGIC_VECTOR(63 downto 0) := (others => '0');
    signal X_L1_PLUS_X_L3, X_L11_PLUS_X_L22, X_L29_PLUS_X_L30, X_L8_PLUS_X_L16, X_L18_PLUS_X_L24 : STD_LOGIC_VECTOR(63 downto 0) := (others => '0');
    signal X_L1_PLUS_X_L3_PLUS_X_L11_PLUS_X_L22, X_L8_PLUS_X_L16_PLUS_X_L18_PLUS_X_L24 : STD_LOGIC_VECTOR(63 downto 0) := (others => '0');
    signal X_L1_PLUS_X_L3_PLUS_X_L11_PLUS_X_L22_PLUS_X_L29_PLUS_X_L30, X_L8_PLUS_X_L16_PLUS_X_L18_PLUS_X_L24_PLUS_X_L26 : STD_LOGIC_VECTOR(63 downto 0) := (others => '0');
    signal X_L1_PLUS_X_L3_PLUS_X_L11_PLUS_X_L22_PLUS_X_L29_PLUS_X_L30_MINUS_X_L8_PLUS_X_L16_PLUS_X_L18_PLUS_X_L24_PLUS_X_L26 : STD_LOGIC_VECTOR(63 downto 0) := (others => '0');
begin
    X_L1  <= "0000000000000000000000000000000" & DIN & "0";
    X_L3  <= "00000000000000000000000000000" & DIN & "000";
    X_L8  <= "000000000000000000000000" & DIN & "00000000";
    X_L11 <= "000000000000000000000" & DIN & "00000000000";
    X_L16 <= "0000000000000000" & DIN & "0000000000000000";
    X_L18 <= "00000000000000" & DIN & "000000000000000000";
    X_L22 <= "0000000000" & DIN & "0000000000000000000000";
    X_L24 <= "00000000" & DIN & "000000000000000000000000";
    X_L26 <= "000000" & DIN & "00000000000000000000000000";
    X_L29 <= "000" & DIN & "00000000000000000000000000000";
    X_L30 <= "00" & DIN & "000000000000000000000000000000";

    X_L1_PLUS_X_L3 <= X_L1 + X_L3;
    X_L11_PLUS_X_L22 <= X_L11 + X_L22;
    X_L29_PLUS_X_L30 <= X_L29 + X_L30;
    X_L8_PLUS_X_L16 <= X_L8 + X_L16;
    X_L18_PLUS_X_L24 <= X_L18 + X_L24;

    X_L1_PLUS_X_L3_PLUS_X_L11_PLUS_X_L22 <= X_L1_PLUS_X_L3 + X_L11_PLUS_X_L22;
    X_L8_PLUS_X_L16_PLUS_X_L18_PLUS_X_L24 <= X_L8_PLUS_X_L16 + X_L18_PLUS_X_L24;

    X_L1_PLUS_X_L3_PLUS_X_L11_PLUS_X_L22_PLUS_X_L29_PLUS_X_L30 <= X_L1_PLUS_X_L3_PLUS_X_L11_PLUS_X_L22 + X_L29_PLUS_X_L30;
    X_L8_PLUS_X_L16_PLUS_X_L18_PLUS_X_L24_PLUS_X_L26 <= X_L8_PLUS_X_L16_PLUS_X_L18_PLUS_X_L24 + X_L26;

    X_L1_PLUS_X_L3_PLUS_X_L11_PLUS_X_L22_PLUS_X_L29_PLUS_X_L30_MINUS_X_L8_PLUS_X_L16_PLUS_X_L18_PLUS_X_L24_PLUS_X_L26 <= X_L1_PLUS_X_L3_PLUS_X_L11_PLUS_X_L22_PLUS_X_L29_PLUS_X_L30 - X_L8_PLUS_X_L16_PLUS_X_L18_PLUS_X_L24_PLUS_X_L26;

    DOUT <= X_L1_PLUS_X_L3_PLUS_X_L11_PLUS_X_L22_PLUS_X_L29_PLUS_X_L30_MINUS_X_L8_PLUS_X_L16_PLUS_X_L18_PLUS_X_L24_PLUS_X_L26(63 downto 32);
end my_mult;
